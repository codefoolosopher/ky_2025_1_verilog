module full_adder (
    input  a,
    input  b,
    input  cin,
    output sum,
    output cout
);
// 코드를 완성 하시오




endmodule
