module half_adder(
	input a,
	input b,
	output sum,
	output carry
);

	// 코드를 완성 하시오



	
endmodule
