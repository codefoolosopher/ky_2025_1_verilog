module tb_full_adder ();

    reg a, b, cin;
    wire sum, cout;

    full_adder dut_FA (
        .a(a),
        .b(b),
        .cin(cin),
        .sum(sum),
        .cout(cout)
    );

    initial begin
        a=0; b=0; cin=0;
        #50 a=1; b=0; cin=0;
        #50 a=0; b=1; cin=0;
        #50 a=1; b=0; cin=0;
        #50 a=1; b=1; cin=0;
        #50 a=0; b=0; cin=1;
        #50 a=1; b=0; cin=1;
        #50 a=0; b=1; cin=1;
        #50 a=1; b=1; cin=1;
        #50 $stop;
    end

endmodule
