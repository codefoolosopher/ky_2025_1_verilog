// exam_dff.v

module dff(  input clk, 
              input din, 
              input rst, 
              output reg q );

//  reg q;
  	// 코드를 완성 하시오




endmodule
