// exam2.v
// verilog calss1 : half_adder circuit
// continuous assignment

`timescale 1ns/10ps

module half_adder2 (
	input a,
	input b,
	output sum,
	output carry
);

	// 코드를 완성 하시오


endmodule
