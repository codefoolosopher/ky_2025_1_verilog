// test bench for half-adder circuit " tb_exam_ha.v "

module tb_ha();

	// 코드를 완성 하시오


endmodule
